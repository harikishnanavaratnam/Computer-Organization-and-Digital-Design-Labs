library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;
-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;
entity Slow_Clk is
Port ( Clk_in : in STD_LOGIC;
 Clk_out : out STD_LOGIC);
end Slow_Clk;
architecture Behavioral of Slow_Clk is
signal count: integer := 1;
signal clk_status: std_logic := '0';
begin
process (Clk_in) begin
if (rising_edge (Clk_in)) then
 count <= count+1;
 if(count = 12) then
 clk_status <= not (clk_status);
 Clk_out <= clk_status;
 count <= 1;
 end if;
end if ;
end process;
end Behavioral;